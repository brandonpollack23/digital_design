library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use ieee.math_real.all;

entity program_counter is
generic
(
	COUNT_WIDTH : natural := log2