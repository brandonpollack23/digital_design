library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std;

entity adder is
  generic (
    WIDTH :     positive := 8);
  port (
    x, y  : in  std_logic_vector(WIDTH-1 downto 0);
    cin   : in  std_logic;
    s     : out std_logic_vector(WIDTH-1 downto 0);
    cout  : out std_logic);
end adder;

architecture RIPPLE_CARRY of adder is

signal carry_vector : std_logic_vector((WIDTH) downto 0);

begin  -- RIPPLE_CARRY
	carry_vector(0) <= cin;
	
	rc_adder : for i in 0 to WIDTH-1 generate
	begin
		ADDER_LSB : if i = 0 generate
		begin
			U0 : entity work.fa port
			map
			(
				a => x(i),
				b => y(i),
				cin => cin,
				cout => carry_vector(i+1),
				sum => s(i)
			);
		end generate ADDER_LSB;
			
		UX : if i > 0 generate
		begin
			UX : entity work.fa port
			map
			(
				a => x(i),
				b => y(i),
				cin => carry_vector(i),
				cout => carry_vector(i+1),
				sum => s(i)
			);
		end generate UX;
	end generate rc_adder;
	
	cout <= carry_vector(WIDTH);
end RIPPLE_CARRY;
		
			


architecture CARRY_LOOKAHEAD of adder is

begin  -- CARRY_LOOKAHEAD

  process(x, y, cin)

    -- generate and propagate bits
    variable g, p : std_logic_vector(WIDTH-1 downto 0);

    -- internal carry bits
    variable carry : std_logic_vector(WIDTH downto 0);

    -- and'd p sequences
    variable p_ands : std_logic_vector(WIDTH-1 downto 0);

  begin

    -- calculate generate (g) and propogate (p) values

    for i in 0 to WIDTH-1 loop
		-- fill in code that defines each g and p bit
		g(i) := x(i) and y(i);

		p(i) := x(i) or y(i);
    end loop;  -- i

    carry(0) := cin;

    -- calculate each carry bit
       
    for i in 1 to WIDTH loop

      -- calculate and'd p terms for ith carry logic      
      -- the index j corresponds to the lowest Pj value in the sequence
      -- e.g., PiPi-1...Pj

      for j in 0 to i-1 loop
        p_ands(j) := '1';

        -- and everything from Pj to Pi-1
        for k in j to i-1 loop
          -- fill code
			p_ands(j) := p_ands(j) and p(k);
			end loop;
      end loop;

      carry(i) := g(i-1);

      -- handle all of the pg minterms
      for j in 1 to i-1 loop
        -- fill in code
		  carry(i) := carry(i) or (g(j-1) and p_ands(j-1));
      end loop;

      -- handle the final propagate of the carry in
      carry(i) := carry(i) or (p_ands(0) and cin);
    end loop;  -- i

    -- set the outputs
    for i in 0 to WIDTH-1 loop
      -- fill in code
		s(i) <= x(i) xor y(i) xor carry(i);
    end loop;  -- i
    
    cout <= carry(WIDTH);

  end process;

end CARRY_LOOKAHEAD;

-- You don't have to change any of the code for the following
-- architecture. However, read the lab instructions to create
-- an RTL schematic of this entity so you can see how the
-- synthesized circuit differs from the previous carry
-- lookahead circuit.

architecture CARRY_LOOKAHEAD_BAD_SYNTHESIS of adder is
begin  -- CARRY_LOOKAHEAD_BAD_SYNTHESIS

  process(x, y, cin)

    -- generate and propagate bits
    variable g, p : std_logic_vector(WIDTH-1 downto 0);

    -- internal carry bits
    variable carry : std_logic_vector(WIDTH downto 0);

  begin

    -- calculate generate (g) and propogate (p) values

    for i in 0 to WIDTH-1 loop
      g(i) := x(i) and y(i);
      p(i) := x(i) or y(i);
    end loop;  -- i

    -- calculate carry bits (the order here is very important)
    -- Problem: defining the carries this way causes the synthesis
    -- tool to chain everything together like a ripple carry.
    -- See RTL view in synthesis tool.
    
    carry(0)     := cin;
    for i in 0 to WIDTH-1 loop
      carry(i+1) := g(i) or (p(i) and carry(i));
    end loop;  -- i

    -- set the outputs

    for i in 0 to WIDTH-1 loop
      s(i) <= x(i) xor y(i) xor carry(i);
    end loop;  -- i

    cout <= carry(WIDTH);

  end process;

end CARRY_LOOKAHEAD_BAD_SYNTHESIS;



architecture HIERARCHICAL of adder is

signal bp0,bp1,bg0,bg1,useless_carry,cout_in_between : std_logic;

begin  -- HIERARCHICAL
	U0 : entity work.cla4 port
	map
	(
		x(3 downto 0) => x(3 downto 0),
		y(3 downto 0) => y(3 downto 0),
		cin => cin,
		cout => useless_carry,
		sum(3 downto 0) => s(3 downto 0),
		bp => bp0,
		bg => bg0
	);
	
	cgen : entity work.cgen2 port
	map
	(
		ci => useless_carry,
		pi => bp0,
		gi => bg0,
		pi_n => bp1,
		gi_n => bg1,
		cout_in_between => cout_in_between,
		cout => cout
	);
	
	U1 : entity work.cla4 port
	map
	(
		x(3 downto 0) => x(7 downto 4),
		y(3 downto 0) => y(7 downto 4),
		cin => cout_in_between,
		sum(3 downto 0) => s(7 downto 4),
		bp => bp1,
		bg => bg1
	);
end HIERARCHICAL;

--architecture extra_credit of adder is
--
--signal bg0,bg1,bp0,bp1,cout_in_between : std_logic;
--
--begin
--	--instantiate two adder_supers and a cgen2, you know what to do
--	--you handsome devil, you
--	ADDER_LOW : entity work.adder_super 
--	generic map
--	(
--		WIDTH => WIDTH/2
--	)
--	port map
--	(
--		x(WIDTH/2-1 downto 0) => x(WIDTH/2-1 downto 0),
--		y(WIDTH/2-1 downto 0) => y(WIDTH/2-1 downto 0),
--		cin => cin,
--		s(WIDTH/2-1 downto 0) => s(WIDTH/2-1 downto 0),
--		bp => bp0,
--		bg => bg0
--	);
--	
--	CGEN : entity work.cgen2
--	port map
--	(
--		ci => cin,
--		pi => bp0,
--		gi => bg0,
--		pi_n => bp1,
--		gi_n => bg1,
--		cout => cout,
--		cout_in_between => cout_in_between
--		--no bp and bg connection on the outside here
--	);
--	
--	ADDER_HIGH : entity work.adder_super
--	generic map
--	(
--		WIDTH => WIDTH/2
--	)
--	port map
--	(
--		x(WIDTH/2-1 downto 0) => x(WIDTH-1 downto WIDTH/2),
--		y(WIDTH/2-1 downto 0) => y(WIDTH-1 downto WIDTH/2),
--		cin => cout_in_between,
--		s(WIDTH/2-1 downto 0) => s(WIDTH-1 downto WIDTH/2),
--		bp => bp1,
--		bg => bg1
--	);
--end extra_credit;